-- PLACEHOLDER, I'M WORKING ON THIS RIGHT NOW
